// DAC handler/interface code for TI TLV5616C digital-analog converter
// Writen by James Dalton 7/6/18

module dac_handler (
    );
    
endmodule